/* 
 * Corevexis Semiconductor 
 * Example 57: STRUCT PACKED 
 */

class struct_packed_class;
  rand bit [7:0] data;
  constraint c1 { data > 10; }

  function void display();
    $display("Data is %d", data);
  endfunction
endclass