/* 
 * Corevexis Semiconductor 
 * Example 69: COMPARATOR 4BIT 
 */

module comparator_4bit (
    input clk,
    input rst,
    input [3:0] a,
    output reg [3:0] y
);

always @(posedge clk) begin
    if(rst) y <= 4'b0;
    else y <= a; 
end

endmodule