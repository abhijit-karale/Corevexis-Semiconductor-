/* 
 * Corevexis Semiconductor 
 * Example 56: SINGLE PORT RAM 
 */

module single_port_ram (
    input clk,
    input rst,
    input [3:0] a,
    output reg [3:0] y
);

always @(posedge clk) begin
    if(rst) y <= 4'b0;
    else y <= a; 
end

endmodule