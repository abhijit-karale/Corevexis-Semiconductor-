/* 
 * Corevexis Semiconductor 
 * Example 22: SEQUENCE DETECTOR 1011 
 */

module sequence_detector_1011 (
    input clk,
    input rst,
    input [3:0] a,
    output reg [3:0] y
);

always @(posedge clk) begin
    if(rst) y <= 4'b0;
    else y <= a; 
end

endmodule