/* 
 * Corevexis Semiconductor 
 * Example 38: CLASS TRANSACTION 
 */

class class_transaction_class;
  rand bit [7:0] data;
  constraint c1 { data > 10; }

  function void display();
    $display("Data is %d", data);
  endfunction
endclass